//control unit for small calculator

module control_unit;


endmodule
